module SWG_design(
  input [9:0] T,
  output [15:0] O
);

  reg [15:0] I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15, I16, I17, I18, I19, I20, I21, I22, I23, I24, I25, I26, I27, I28, I29, I30, I31, I32, I33, I34, I35, I36, I37, I38, I39, I40, I41, I42, I43, I44, I45, I46, I47, I48, I49, I50, I51, I52, I53, I54, I55, I56, I57, I58, I59, I60, I61, I62, I63;

  MUX16_64_design m1(
    .I0(I0), .I1(I1), .I2(I2), .I3(I3), .I4(I4), .I5(I5), .I6(I6), .I7(I7), .I8(I8), .I9(I9), .I10(I10), .I11(I11), .I12(I12), .I13(I13), .I14(I14), .I15(I15),
    .I16(I16), .I17(I17), .I18(I18), .I19(I19), .I20(I20), .I21(I21), .I22(I22), .I23(I23), .I24(I24), .I25(I25), .I26(I26), .I27(I27), .I28(I28), .I29(I29), .I30(I30), .I31(I31),
    .I32(I32), .I33(I33), .I34(I34), .I35(I35), .I36(I36), .I37(I37), .I38(I38), .I39(I39), .I40(I40), .I41(I41), .I42(I42), .I43(I43), .I44(I44), .I45(I45), .I46(I46), .I47(I47),
    .I48(I48), .I49(I49), .I50(I50), .I51(I51), .I52(I52), .I53(I53), .I54(I54), .I55(I55), .I56(I56), .I57(I57), .I58(I58), .I59(I59), .I60(I60), .I61(I61), .I62(I62), .I63(I63),
    .T(T), .O(O)
  );

  initial begin
    I0  = 1000; I1  = 1098; I2  = 1195; I3  = 1290;
    I4  = 1383; I5  = 1471; I6  = 1556; I7  = 1634;
    I8  = 1707; I9  = 1773; I10 = 1831; I11 = 1882;
    I12 = 1924; I13 = 1957; I14 = 1981; I15 = 1995;
    I16 = 2000; I17 = 1995; I18 = 1981; I19 = 1957;
    I20 = 1924; I21 = 1882; I22 = 1831; I23 = 1773;
    I24 = 1707; I25 = 1634; I26 = 1556; I27 = 1471;
    I28 = 1383; I29 = 1290; I30 = 1195; I31 = 1098; 
    I32 = 1000; I33 = 902;  I34 = 805;  I35 = 710; 
    I36 = 617;  I37 = 529;  I38 = 444;  I39 = 366; 
    I40 = 293;  I41 = 227;  I42 = 169;  I43 = 118; 
    I44 = 76;   I45 = 43;   I46 = 19;   I47 = 5;
    I48 = 0;    I49 = 5;    I50 = 19;   I51 = 43; 
    I52 = 76;   I53 = 118;  I54 = 169;  I55 = 227; 
    I56 = 293;  I57 = 366;  I58 = 444;  I59 = 529; 
    I60 = 617;  I61 = 710;  I62 = 805;  I63 = 902;
  end

endmodule
