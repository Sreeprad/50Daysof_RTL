module FA_TB;

    reg A, B, C;

    wire Sum, Carry;
    
    FA_design uut(A, B, C, Sum, Carry);

    initial begin
        A = 0; B = 0; C = 0; #10;
        A = 0; B = 1; C = 0; #10;
        A = 1; B = 0; C = 0; #10;
        A = 1; B = 1; C = 0; #10;
        A = 0; B = 0; C = 1; #10;
        A = 0; B = 1; C = 1; #10;
        A = 1; B = 0; C = 1; #10;
        A = 1; B = 1; C = 1; #10;
        $finish();
    end

endmodule
